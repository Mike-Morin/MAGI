.title KiCad schematic
R1 +9V Net-_C1-Pad2_ 10K
R2 Net-_C1-Pad2_ -9V 10K
C1 +9V Net-_C1-Pad2_ 10u
C2 Net-_C1-Pad2_ -9V 10u
U1 Net-_C4-Pad2_ GND Net-_C1-Pad2_ -9V GND Net-_U1-Pad6_ Net-_U1-Pad6_ +9V NE5532
U2 Net-_R3-Pad2_ Net-_C4-Pad1_ Net-_C4-Pad1_ +9V NC_01 Net-_C4-Pad1_ Net-_C4-Pad1_ NC_02 LM334
Q1 Net-_C4-Pad2_ Net-_Q1-Pad2_ Net-_C4-Pad1_ 2N2222
R5 Net-_C4-Pad1_ Net-_Q1-Pad2_ 1.1K
RV1 Net-_Q1-Pad2_ Net-_C4-Pad2_ Net-_C4-Pad2_ 1K
R4 Net-_C4-Pad2_ -9V 5.6K
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ 10n
Q2 Net-_C4-Pad1_ +9V Net-_Q2-Pad3_ TIP122
Q3 Net-_C4-Pad2_ Net-_Q3-Pad2_ -9V TIP127
R6 Net-_Q2-Pad3_ GND 1R
R7 GND Net-_Q3-Pad2_ 1R
C5 +9V GND 220u
C6 GND -9V 220u
R3 +9V Net-_R3-Pad2_ 14R
C3 +9V -9V 100n
J2 +9V GND -9V Power_Header
J1 -9V +9V Conn_01x02
.end
